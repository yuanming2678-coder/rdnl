.global VSS VDD

.subckt ALU4 A0 A1 A2 A3 B0 B1 B2 B3 M0 M1 S0 S1 S2 S3 COUT
XAND0 A0 B0 AND0 AND2
XAND1 A1 B1 AND1 AND2
XAND2 A2 B2 AND2 AND2
XAND3 A3 B3 AND3 AND2
XFA0 A0 BB0 M0 SUM0 C0 FULLADDER
XFA1 A1 BB1 C0 SUM1 C1 FULLADDER
XFA2 A2 BB2 C1 SUM2 C2 FULLADDER
XFA3 A3 BB3 C2 SUM3 COUT FULLADDER
XM0A SUM0 AND0 M1 S0 MUX2
XM0B S0 OR0 M0 S0 MUX2
XM1A SUM1 AND1 M1 S1 MUX2
XM1B S1 OR1 M0 S1 MUX2
XM2A SUM2 AND2 M1 S2 MUX2
XM2B S2 OR2 M0 S2 MUX2
XM3A SUM3 AND3 M1 S3 MUX2
XM3B S3 OR3 M0 S3 MUX2
XMUX0 B0 NB0 M1 BB0 MUX2
XMUX1 B1 NB1 M1 BB1 MUX2
XMUX2 B2 NB2 M1 BB2 MUX2
XMUX3 B3 NB3 M1 BB3 MUX2
XNOT0 B0 NB0 NOT
XNOT1 B1 NB1 NOT
XNOT2 B2 NB2 NOT
XNOT3 B3 NB3 NOT
XOR0 A0 B0 XOR0 XOR2
XOR1 XOR0 B0 OR0 OR2
XOR2 A1 B1 XOR1 XOR2
XOR3 XOR1 B1 OR1 OR2
XOR4 A2 B2 XOR2 XOR2
XOR5 XOR2 B2 OR2 OR2
XOR6 A3 B3 XOR3 XOR2
XOR7 XOR3 B3 OR3 OR2
.ends ALU4

.subckt AND2 A B Y
M1 N1 A VSS VSS NMOS W=1u L=0.18u
M2 Y B N1 VSS NMOS W=1u L=0.18u
M3 Y A VDD VDD PMOS W=2u L=0.18u
M4 Y B VDD VDD PMOS W=2u L=0.18u
.ends AND2

.subckt FULLADDER A B CIN SUM COUT
X1 A B S1 XOR2
X2 S1 CIN SUM XOR2
X3 A B T1 AND2
X4 B CIN T2 AND2
X5 A CIN T3 AND2
X6 T1 T2 T4 OR2
X7 T4 T3 COUT OR2
.ends FULLADDER

.subckt MUX2 A B SEL Y
X1 SEL NSEL NOT
X2 A NSEL T1 AND2
X3 B SEL T2 AND2
X4 T1 T2 Y OR2
.ends MUX2

.subckt NAND2 A B Y
M1 Y A VSS VSS NMOS W=1u L=0.18u
M2 Y B VSS VSS NMOS W=1u L=0.18u
M3 Y A VDD VDD PMOS W=2u L=0.18u
M4 Y B VDD VDD PMOS W=2u L=0.18u
.ends NAND2

.subckt NOT A Y
M1 Y A VSS VSS NMOS W=1u L=0.18u
M2 Y A VDD VDD PMOS W=2u L=0.18u
.ends NOT

.subckt OR2 A B Y
M1 Y A VSS VSS NMOS W=1u L=0.18u
M2 Y B VSS VSS NMOS W=1u L=0.18u
M3 N1 A VDD VDD PMOS W=2u L=0.18u
M4 Y B N1 VDD PMOS W=2u L=0.18u
.ends OR2

.subckt XOR2 A B Y
X1 A B T1 NAND2
X2 A T1 T2 NAND2
X3 B T1 T3 NAND2
X4 T2 T3 Y NAND2
.ends XOR2

cs0 s0 VSS 1f
ra0 a0 VSS 1k
rb1 a1 VSS 1k
vvdd VDD VSS 2.2
vvdd VSS 0 0
xalu4 a0 a1 a2 a3 b0 b1 b2 b3 mode[0] mode[1] s0 s1 s2 s3 cout ALU4
